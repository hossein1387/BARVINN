../../../pito_riscv/verification/lib/utils/pito_pkg.sv