../../../pito_riscv/verification/lib/utils/rv32_utils.sv